module scope(
	
);

endmodule // scope
